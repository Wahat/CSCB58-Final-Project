// mux module winner
// 1 for winner
// 0 for loser
// input: switch, output to hex

module endgame (reg_win, reg_lose, in, out, out2);
  input in;
  output [6:0] win;
  output [6:0] lose;

  m =



endmodule;
