// Draw black square over play area to reset
module clearscreen(in, out);
  input in;
  output out;

endmodule
